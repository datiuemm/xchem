** sch_path: /home/datdt/xchem/xchem/inverter.sch
.subckt inverter VDD A Y VSS
*.PININFO A:I VDD:B VSS:B Y:O
M1 Y A VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
M2 Y A VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends
.end
