** sch_path: /home/datdt/xchem/xchem/Bai1_Basic_RLC.sch
**.subckt Bai1_Basic_RLC
C1 A B 50nF m=1
R1 A 0 1k m=1
E1 C 0 VOL=' 3*cos(time*time*time*1e11) '
L1 B C 10mH m=1
**** begin user architecture code

.tran 10n 2000u uic
.save all

**** end user architecture code
**.ends
.end
